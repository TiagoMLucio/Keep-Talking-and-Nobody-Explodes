library ieee;
use ieee.std_logic_1164.all;

entity circuito_jogo_base is
    port (
        clock       : in std_logic;
        reset       : in std_logic;
        iniciar     : in std_logic;
        botoes      : in std_logic_vector (3 downto 0);
        leds        : out std_logic_vector (3 downto 0);
        pronto      : out std_logic;
        ganhou      : out std_logic;
        perdeu      : out std_logic;
        db_clock    : out std_logic;
        db_igual    : out std_logic;
        db_timeout  : out std_logic;
        db_contagem : out std_logic_vector (6 downto 0);
        db_memoria  : out std_logic_vector (6 downto 0);
        db_jogada   : out std_logic_vector (6 downto 0);
        db_rodada   : out std_logic_vector (6 downto 0);
        db_estado   : out std_logic_vector (6 downto 0)
    );
end entity;
architecture estrutural of circuito_jogo_base is

    signal zeraE, zeraCR, zeraT, contaE, contaCR, contaT, escreve, limpaRC, registraRC, jogada_correta, enderecoIgualRodada, fimE, fimL, fimT, jogada_feita : std_logic;
    signal db_contagem_t, db_jogada_t, db_rodada_t, db_estado_t, memoria_s                                                                                  : std_logic_vector (3 downto 0);

    component fluxo_dados
        port (
            clock               : in std_logic;
            zeraE               : in std_logic;
            zeraCR              : in std_logic;
            zeraT               : in std_logic;
            contaE              : in std_logic;
            contaCR             : in std_logic;
            contaT              : in std_logic;
            escreve             : in std_logic;
            limpaRC             : in std_logic;
            registraRC          : in std_logic;
            chaves              : in std_logic_vector (3 downto 0);
            jogada_correta      : out std_logic;
            enderecoIgualRodada : out std_logic;
            fimE                : out std_logic;
            fimL                : out std_logic;
            fimT                : out std_logic;
            jogada_feita        : out std_logic;
            memoria_s           : out std_logic_vector (3 downto 0);
            db_contagem         : out std_logic_vector (3 downto 0);
            db_rodada           : out std_logic_vector (3 downto 0);
            db_jogada           : out std_logic_vector (3 downto 0)
        );
    end component;

    component unidade_controle is
        port (
            clock               : in std_logic;
            reset               : in std_logic;
            iniciar             : in std_logic;
            fimL                : in std_logic;
            fimT                : in std_logic;
            jogada_feita        : in std_logic;
            enderecoIgualRodada : in std_logic;
            jogada_correta      : in std_logic;
            contaE              : out std_logic;
            contaT              : out std_logic;
            contaCR             : out std_logic;
            registraRC          : out std_logic;
            zeraE               : out std_logic;
            zeraT               : out std_logic;
            zeraCR              : out std_logic;
            limpaRC             : out std_logic;
            pronto              : out std_logic;
            ganhou              : out std_logic;
            perdeu              : out std_logic;
            db_timeout          : out std_logic;
            db_estado           : out std_logic_vector(3 downto 0)
        );
    end component;

    component hexa7seg is
        port (
            hexa : in std_logic_vector(3 downto 0);
            sseg : out std_logic_vector(6 downto 0)
        );
    end component;

begin

    fd : fluxo_dados
    port map(
        clock               => clock,
        zeraE               => zeraE,
        zeraCR              => zeraCR,
        zeraT               => zeraT,
        contaE              => contaE,
        contaCR             => contaCR,
        contaT              => contaT,
        escreve             => escreve,
        limpaRC             => limpaRC,
        registraRC          => registraRC,
        chaves              => botoes,
        jogada_correta      => jogada_correta,
        enderecoIgualRodada => enderecoIgualRodada,
        fimE                => fimE,
        fimL                => fimL,
        fimT                => fimT,
        jogada_feita        => jogada_feita,
        memoria_s           => memoria_s,
        db_contagem         => db_contagem_t,
        db_rodada           => db_rodada_t,
        db_jogada           => db_jogada_t
    );

    uc : unidade_controle
    port map(
        clock               => clock,
        reset               => reset,
        iniciar             => iniciar,
        fimL                => fimL,
        fimT                => fimT,
        jogada_feita        => jogada_feita,
        enderecoIgualRodada => enderecoIgualRodada,
        jogada_correta      => jogada_correta,
        contaE              => contaE,
        contaT              => contaT,
        contaCR             => contaCR,
        registraRC          => registraRC,
        zeraE               => zeraE,
        zeraT               => zeraT,
        zeraCR              => zeraCR,
        limpaRC             => limpaRC,
        pronto              => pronto,
        ganhou              => ganhou,
        perdeu              => perdeu,
        db_timeout          => db_timeout,
        db_estado           => db_estado_t
    );

    HEX0 : hexa7seg
    port map(
        hexa => db_contagem_t,
        sseg => db_contagem
    );

    HEX1 : hexa7seg
    port map(
        hexa => memoria_s,
        sseg => db_memoria
    );

    HEX2 : hexa7seg
    port map(
        hexa => db_jogada_t,
        sseg => db_jogada
    );

    HEX3 : hexa7seg
    port map(
        hexa => db_rodada_t,
        sseg => db_rodada
    );

    HEX5 : hexa7seg
    port map(
        hexa => db_estado_t,
        sseg => db_estado
    );

    db_igual <= jogada_correta;
    db_clock <= clock;

end architecture estrutural;
